`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 08/18/2022 07:37:56 PM
// Design Name: 
// Module Name: module_memoria
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module module_memoria_spi(
    input   logic                           clk_i,
    input   logic                           rst_i,
    input   logic                           we_i,
    input  pkg_global:: bitsh_t             addr_rs1_i,
    input  pkg_global:: bitsh_t             addr_rd_i,
    input  pkg_global:: bits_width          data_in_i,
    output pkg_global:: bits_width          rs1_o
                     );
    
    import                                  pkg_global::*;
    
    
    logic [63 : 0][31 : 0]                 memoria;
    
    always @ ( posedge clk_i ) begin
     if   ( rst_i )  memoria <=          '0;
     else begin 
            if ( we_i ) begin
                memoria [ addr_rd_i ] <= data_in_i; 
            end
     end
    end
    
    //Logica de salida
    always_comb begin
        rs1_o = memoria [ addr_rs1_i ];
    end
endmodule
